module de0_nano_toplevel (
    input        user_50mhz_clk, // CLOCK_50 [PIN_R8]
    input        user_rst_n, // Key 0 [PIN_J15]
       
    input        user_button_n, // key 1 [PIN_E1]
    input  [3:0] dip_switches,  // Active DOWN/ON [PIN_M15, PIN_B9, PIN_T8, PIN_M1]

    output [7:0] green_leds, // [PIN_L3, PIN_B1, PIN_F3, PIN_D1, PIN_A11, PIN_B13, PIN_A13, PIN_A15]

    output       sclk, // ADC_SCLK [PIN_B14]
    output       cs_n, // ADC_CS_N [PIN_A10]
    output       copi, // ADC_SADDR [PIN_B10]
    input        cipo  // ADC_SDAT [PIN_A9]

    //TODO: Finish I2C Controller to use with the ADXL345
    // // ADXL345 Accelerometer
    // output       i2c_sclk,
    // inout        i2c_sdat,
    // input        accel_interrupt
);

//? System Control
    //                                                                       //
    //* Common Connections and Parameters
        localparam integer Reset_Pulse_Length = 8;
        localparam integer Reset_Delay_Cycles = 1024; // How many cycles after a reset is detected, is it actually forwarded to the rest of the system.
        localparam integer Button_Validation_Wait_Cycles = 2_500_000; // 50ms @ 50Mhz
        localparam integer Button_Lockout_Cycles = 5_000_000; // 100ms of a second @ 50Mhz
    
    // These are connections that are used either before they are driven in this section, or connect to something outside this module
        wire power_on_reset_n;
        
        wire async_rst;
        wire clk_lock;

        wire clk_sys;
        wire clk_en_sys;
        wire sync_rst_sys;
        wire init_sys;
    //                                                                       //
    //* Power-On-Reset Detection
    //! Note: This will be FPGA-Specific and will need to be generated by a chips respective tooling suite.
    /*
    On a Cyclone IV or V, you can use the following to detect a power-up. This
    works as the default configuration for both generations trigger a localized
    async_clear for every register
    */
        reg  [3:0] power_on_reset_vector_current;
        wire       por_saturation_check = power_on_reset_vector_current == 4'hF;
        wire       power_on_reset_lsb = power_on_reset_vector_current[0] || ~por_saturation_check;
        wire [3:0] power_on_reset_vector_next = {power_on_reset_vector_current[2:0], power_on_reset_lsb};
        always_ff @(posedge user_50mhz_clk) begin
            power_on_reset_vector_current <= power_on_reset_vector_next;
        end
        assign power_on_reset_n = ~power_on_reset_vector_current[3];
    //                                                                       //
    //* Reset Synchronization + Power-On-Reset Detection
        reset_control #(
            .Reset_Pulse_Length          (Reset_Pulse_Length),
            .Reset_Delay_Cycles          (Reset_Delay_Cycles),
            .Press_Validation_Wait_Cycles(Button_Validation_Wait_Cycles),
            .Release_Lockout_Cycles      (Button_Lockout_Cycles)
        ) reset_controller (
            .user_clk  (user_50mhz_clk),
            .user_rst_n(user_rst_n),
            .por_n     (power_on_reset_n),
            .async_rst (async_rst)
        );
    //                                                                       //
    //* PLL - Clock Control
    // input_clk    - 50Mhz
    // sys_clk (c0) - 50Mhz
        pll clock_generation (
    	    .areset(async_rst),
    	    .inclk0(user_50mhz_clk),
    	    .c0    (clk_sys),
    	    .locked(clk_lock)
        );
    //                                                                       //
    //* Sys Clock Domain Control
        domain_control sys_domain_control (
            .clk          (clk_sys),
            .async_rst    (async_rst),
            .domain_enable(clk_lock),
            .clk_en       (clk_en_sys),
            .sync_rst     (sync_rst_sys),
            .init         (init_sys)
        );
    //                                                                       //
//?

//? IO Drivers
    //                                                                       //
    //* Common Connections
        localparam integer Pulse_Length = 1;
        localparam integer Repeat_Wait_Cycles = 10_000_000; // 250ms of a second @ 50Mhz

        wire       button_pulse;
        wire [3:0] switch_states;
        wire [7:0] led_states;

        wire update_ack;

        wire [7:0][11:0] adc_channels_data;
        wire       [7:0] adc_channels_valid;

        wire copi_d;
        wire copi_en;

    //                                                                       //
    //* Button
        monostable_debouncer #(
            .Press_Validation_Wait_Cycles(Button_Validation_Wait_Cycles),
            .Release_Lockout_Cycles      (Button_Lockout_Cycles),
            .Pulse_Length                (Pulse_Length),
            .Repeat_Wait_Cycles          (Repeat_Wait_Cycles)
        ) user_button_control (
            .clk            (clk_sys),
            .clk_en         (clk_en_sys),
            .sync_rst       (sync_rst_sys),
            .repeat_en      (1'b1),
            .io_in          (~user_button_n),
            .debounced_pulse(button_pulse)
        );
    //                                                                       //
    //* Dip Switches
        de0_nano_dip_switches #(
            .Validation_Wait_Cycles(Button_Validation_Wait_Cycles),
            .Lockout_Cycles        (Button_Lockout_Cycles)
        ) dip_switche_control (
            .clk         (clk_sys),
            .clk_en      (clk_en_sys),
            .sync_rst    (sync_rst_sys),
            .dip_switches(dip_switches),
            .state_out   (switch_states)
        );
    //                                                                       //
    //* Green LEDs
        logic  [7:0] selected_led_source;
        always_comb begin : selected_led_source_mux
            case (switch_states)
                4'h0   : selected_led_source = adc_channels_data[0][7:0];
                4'h1   : selected_led_source = adc_channels_data[1][7:0];
                4'h2   : selected_led_source = adc_channels_data[2][7:0];
                4'h3   : selected_led_source = adc_channels_data[3][7:0];
                4'h4   : selected_led_source = adc_channels_data[4][7:0];
                4'h5   : selected_led_source = adc_channels_data[5][7:0];
                4'h6   : selected_led_source = adc_channels_data[6][7:0];
                4'h7   : selected_led_source = adc_channels_data[7][7:0];
                4'h8   : selected_led_source = {adc_channels_valid[0], 3'd0, adc_channels_data[0][11:8]};
                4'h9   : selected_led_source = {adc_channels_valid[1], 3'd0, adc_channels_data[1][11:8]};
                4'hA   : selected_led_source = {adc_channels_valid[2], 3'd0, adc_channels_data[2][11:8]};
                4'hB   : selected_led_source = {adc_channels_valid[3], 3'd0, adc_channels_data[3][11:8]};
                4'hC   : selected_led_source = {adc_channels_valid[4], 3'd0, adc_channels_data[4][11:8]};
                4'hD   : selected_led_source = {adc_channels_valid[5], 3'd0, adc_channels_data[5][11:8]};
                4'hE   : selected_led_source = {adc_channels_valid[6], 3'd0, adc_channels_data[6][11:8]};
                4'hF   : selected_led_source = {adc_channels_valid[7], 3'd0, adc_channels_data[7][11:8]};
                default: selected_led_source = 8'd0;
            endcase
        end

        de0_nano_leds_top_generic led_controller (
            .clk        (clk_sys),
            .clk_en     (clk_en_sys),
            .sync_rst   (sync_rst_sys),
            .data_in    (selected_led_source),
            .update_leds(1'b1),
            .leds_out   (green_leds)
        );
    //                                                                       //
    //* Analog to Digital Converter
        wire single_update_req = ~switch_states[3] && button_pulse;
        wire burst_update_req = switch_states[3] && button_pulse;

        reg  [2:0] adc_channel_current;
        wire [2:0] adc_channel_next = sync_rst_sys ? 3'd0 : (adc_channel_current + 3'd1);
        wire        adc_channel_trigger = sync_rst_sys || (clk_en_sys && single_update_req && update_ack);
        always_ff @(posedge clk_sys) begin
            if (adc_channel_trigger) begin
                adc_channel_current <= adc_channel_next;
            end
        end
        
        adc128s022_top_generic adc_controller (
            .clk              (clk_sys),
            .clk_en           (clk_en_sys),
            .sync_rst         (sync_rst_sys),
            .single_update_req(single_update_req),
            .burst_update_req (burst_update_req),
            .update_ack       (update_ack),
            .channel_addr     (adc_channel_current),
            .channels_out     (adc_channels_data),
            .channel_valid    (adc_channels_valid),
            .sclk             (sclk),
            .cs_n             (cs_n),
            .copi             (copi_d),
            .copi_en          (copi_en),
            .cipo             (cipo)
        );

        io_out_buf_iobuf_out_d5t ( 
        	.datain (copi_d),
        	.dataout(copi_en),
        	.oe     (copi)
        );
    //                                                                       //
//?

//? Platform Independent

//?

endmodule : de0_nano_toplevel
