module de10_standard_toplevel (
    input        user_50mhz_clk,
    input        user_rst_n, // Key 0 [PIN_AJ4]
       
    input  [2:0] user_buttons_n, // key 3:1 [PIN_AA15, PIN_AA14, PIN_AK4]
    
);

// TODO: Still need to add example code to this.

//? System Control
    //                                                                       //
    //* Common Connections and Parameters
        localparam integer Reset_Pulse_Length = 8;
        localparam integer Reset_Delay_Cycles = 1024; // How many cycles after a reset is detected, is it actually forwarded to the rest of the system.
        localparam integer Press_Validation_Wait_Cycles = 3_500; // 1ms @ 35Mhz
        localparam integer Release_Lockout_Cycles = 350_000; // 1/10th of a second @ 35Mhz
    
    // These are connections that are used either before they are driven in this section, or connect to something outside this module
        wire power_on_reset_n;
        
        wire async_rst;
        wire clk_lock;

        wire clk_sys;
        wire clk_en_sys;
        wire sync_rst_sys;
        wire init_sys;
    //                                                                       //
    //* Power-On-Reset Detection
    //! Note: This will be FPGA-Specific and will need to be generated by a chips respective tooling suite.
    /*
    On a Cyclone IV or V, you can use the following to detect a power-up. This
    works as the default configuration for both generations trigger a localized
    async_clear for every register
    */
        reg  [3:0] power_on_reset_vector_current;
        wire       por_saturation_check = power_on_reset_vector_current == 4'hF;
        wire       power_on_reset_lsb = power_on_reset_vector_current[0] || ~por_saturation_check;
        wire [3:0] power_on_reset_vector_next = {power_on_reset_vector_current[2:0], power_on_reset_lsb};
        always_ff @(posedge user_50mhz_clk) begin
            power_on_reset_vector_current <= power_on_reset_vector_next;
        end
        assign power_on_reset_n = ~power_on_reset_vector_current[3];
    //                                                                       //
    //* Reset Synchronization + Power-On-Reset Detection
        reset_control #(
            .Reset_Pulse_Length          (Reset_Pulse_Length),
            .Reset_Delay_Cycles          (Reset_Delay_Cycles),
            .Press_Validation_Wait_Cycles(Press_Validation_Wait_Cycles),
            .Release_Lockout_Cycles      (Release_Lockout_Cycles)
        ) reset_controller (
            .user_clk  (user_50mhz_clk),
            .user_rst_n(user_rst_n),
            .por_n     (power_on_reset_n),
            .async_rst (async_rst)
        );
    //                                                                       //
    //* PLL - Clock Control
    // input_clk    - 50Mhz
    // sys_clk (c0) - 35Mhz
        pll clock_generation (
    	    .rst     (async_rst),
    	    .refclk  (user_50mhz_clk),
    	    .outclk_0(clk_sys),
    	    .locked  (clk_lock)
        );
    //                                                                       //
    //* Sys Clock Domain Control
        domain_control sys_domain_control (
            .clk          (clk_sys),
            .async_rst    (async_rst),
            .domain_enable(clk_lock),
            .clk_en       (clk_en_sys),
            .sync_rst     (sync_rst_sys),
            .init         (init_sys)
        );
    //                                                                       //
//?

//? IO Drivers
    //                                                                       //

    //                                                                       //
//?

//? Platform Independent

//?

endmodule : de10_standard_toplevel
