/**
 *  Module: platform_independent_top_generic
 *
 *  About: Use this to put any code that you want to run on different target FPGAs/Boards.
 *
**/
module platform_independent_top_generic (
    // 25Mhz Clock
    input        clk_sys,
    input        clk_en_sys,
    input        sync_rst_sys,
    input        init_sys

);












endmodule : platform_independent_top_generic
