module cyclone_v_gx_toplevel (
    input        user_50mhz_clk,
    input        user_rst_n,
       
    input  [3:0] user_buttons_n,
    output [2:0] green_leds,
    output [6:0] hex_0,
    output [6:0] hex_1,
    output [6:0] hex_2,
    output [6:0] hex_3
);

//? System Control
    //                                                                       //
    //* Common Connections and Parameters
        localparam integer Reset_Pulse_Length = 8;
        localparam integer Reset_Delay_Cycles = 1024; // How many cycles after a reset is detected, is it actually forwarded to the rest of the system.
        localparam integer Press_Validation_Wait_Cycles = 3_500; // 1ms @ 35Mhz
        localparam integer Release_Lockout_Cycles = 350_000; // 1/10th of a second @ 35Mhz
    
    // These are connections that are used either before they are driven in this section, or connect to something outside this module
        wire power_on_reset_n;
        
        wire async_rst;
        wire clk_lock;

        wire clk_sys;
        wire clk_en_sys;
        wire sync_rst_sys;
        wire init_sys;
    //                                                                       //
    //* Power-On-Reset Detection
    //! Note: This will be FPGA-Specific and will need to be generated by a chips respective tooling suite.
    /*
    On a Cyclone IV or V, you can use the following to detect a power-up. This
    works as the default configuration for both generations trigger a localized
    async_clear for every register
    */
        reg  [3:0] power_on_reset_vector_current;
        wire       por_saturation_check = power_on_reset_vector_current == 4'hF;
        wire       power_on_reset_lsb = power_on_reset_vector_current[0] || ~por_saturation_check;
        wire [3:0] power_on_reset_vector_next = {power_on_reset_vector_current[2:0], power_on_reset_lsb};
        always_ff @(posedge user_50mhz_clk) begin
            power_on_reset_vector_current <= power_on_reset_vector_next;
        end
        assign power_on_reset_n = ~power_on_reset_vector_current[3];
    //                                                                       //
    //* Reset Synchronization + Power-On-Reset Detection
        reset_control #(
            .Reset_Pulse_Length          (Reset_Pulse_Length),
            .Reset_Delay_Cycles          (Reset_Delay_Cycles),
            .Press_Validation_Wait_Cycles(Press_Validation_Wait_Cycles),
            .Release_Lockout_Cycles      (Release_Lockout_Cycles)
        ) reset_controller (
            .user_clk      (user_50mhz_clk),
            .user_rst_n    (user_rst_n),
            .por_n         (power_on_reset_n),
            .async_rst     (async_rst)
        );
    //                                                                       //
    //* PLL - Clock Control
    // input_clk    - 50Mhz
    // sys_clk (c0) - 35Mhz
        pll clock_generation (
    	    .rst     (async_rst),
    	    .refclk  (user_50mhz_clk),
    	    .outclk_0(clk_sys),
    	    .locked  (clk_lock)
        );
    //                                                                       //
    //* Sys Clock Domain Control
        domain_control sys_domain_control (
            .clk          (clk_sys),
            .async_rst    (async_rst),
            .domain_enable(clk_lock),
            .clk_en       (clk_en_sys),
            .sync_rst     (sync_rst_sys),
            .init         (init_sys)
        );
    //                                                                       //
//?

//? IO Drivers
    //                                                                       //
    //* Common Connections
        wire [3:0] button_pulse_vector; // {Up(Inc), Down(Dec), Right(Invert LED), Sel(Clear)}

        wire [2:0] count_lower;
        wire [6:0] digit_3;   
    //                                                                       //
    //* Buttons
        buttons_top_generic dpad_debouncing (
            .clk                (clk_sys),
            .clk_en             (clk_en_sys),
            .sync_rst           (sync_rst_sys),
            .buttons_n          (user_buttons_n),
            .button_pulse_vector(button_pulse_vector)
        );
    //                                                                       //
    //* Green LED Test
    //TODO: Update this to test *ALL* LEDs
        rgb_test_top_generic rgb_driver (
            .clk             (clk_sys),
            .clk_en          (clk_en_sys),
            .sync_rst        (sync_rst_sys),
            .count_lower     (count_lower),
            .invert_led_state(button_pulse_vector[0]),
            .digit_3         (digit_3),
            .rgb_state       (green_leds)
        );
    //                                                                       //
    //* Seven Segments
        seven_segment_top_generic seven_segment_driver (
            .clk         (clk_sys),
            .clk_en      (clk_en_sys),
            .sync_rst    (sync_rst_sys),
            .clk_pps     (32'd25_000_000),
            .increment   (button_pulse_vector[3]),
            .decrement   (button_pulse_vector[2]),
            .clear       (button_pulse_vector[1]),
            .count_lower (count_lower),
            .digit_3_in  (digit_3),
            .digit_0     (hex_0),
            .digit_1     (hex_1),
            .digit_2     (hex_2),
            .digit_3     (hex_3),
            .segments    (), //! Not used for Cyclone V GX Starter Kit
            .digit_select()  //! Not used for Cyclone V GX Starter Kit
        );
    //                                                                       //
//?

//? Platform Independent

//?

endmodule : cyclone_v_gx_toplevel
